package switch_pkg;
    `include "./switch_item.sv"
    `include "./generator.sv"
  
    `include "./driver.sv"
    `include "./monitor.sv"

    `include "./scoreboard.sv"
    `include "./env.sv"
    `include "./test.sv"
endpackage